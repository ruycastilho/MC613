LIBRARY ieee ; 
USE ieee.std_logic_1164.all;

ENTITY ex1 IS 
	PORT (m:		IN STD_LOGIC;
			n:		IN STD_LOGIC;
			A:		IN STD_LOGIC;
			B:		IN STD_LOGIC;
			clk:	IN STD_LOGIC;
			Q1: 	OUT STD_LOGIC;
			Q2: 	OUT STD_LOGIC;
			Q3: 	OUT STD_LOGIC;
			Q4: 	OUT STD_LOGIC;
			Q5: 	OUT STD_LOGIC;
			Q6: 	OUT STD_LOGIC);
END ex1;

ARCHITECTURE Behavior OF ex1 IS
	BEGIN

				
END Behavior ;